class axi_vip_cfg extends uvm_object;
  `uvm_object_utils(axi_vip_cfg)
  
  
  
  function new(string name ="");
    super.new(name);
  endfunction
  
  
endclass