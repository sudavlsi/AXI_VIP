`include "tests/axi_vip_base_test.sv"
